// Mandatory file to be able to launch SVUT flow
`include "svut_h.sv"

// Specify here the module to load or setup the path in files.f
`include "Adder.v"

`timescale 1 ns / 1 ps

module Adder_unit_test_KO;

    `SVUT_SETUP

    parameter WIDTH = 8;

    reg             aclk;
    reg             arstn;
    reg             clr;
    reg             inc;
    reg [WIDTH-1:0] out;

    Adder
    #(
    WIDTH
    )
    dut
    (
    aclk,
    arstn,
    clr,
    inc,
    out
    );

    // An example to create a clock
    initial aclk = 0;
    always #2 aclk <= ~aclk;

    // An example to dump data for visualization
    initial $dumpvars(0, Adder_unit_test_KO);

    task setup();
    begin
        // setup() runs when a test begins
        inc = 1'b0;
        clr = 1'b0;
        arstn = 1'b0;
        #100;
        arstn = 1'b1;
    end
    endtask

    task teardown();
    begin
        // teardown() runs when a test ends
    end
    endtask

    `TEST_SUITE("")

        /* Available macros:

               - `INFO("message"); Print a grey message
               - `SUCCESS("message"); Print a green message
               - `WARNING("message"); Print an orange message and increment warning counter
               - `CRITICAL("message"); Print an pink message and increment critical counter
               - `ERROR("message"); Print a red message and increment error counter
               - `FAIL_IF(aSignal); Increment error counter if evaluaton is positive
               - `FAIL_IF_NOT(aSignal); Increment error coutner if evaluation is false
               - `FAIL_IF_EQUAL(aSignal, 23); Increment error counter if evaluation is equal
               - `FAIL_IF_NOT_EQUAL(aSignal, 45); Increment error counter if evaluation is not equal
        */

        /* Available flag:

               - `LAST_STATUS: tied to 1 is last macros has been asserted, else tied to 0
        */

    `UNIT_TEST("REGRESSION")

        `INFO("Start REGRESSION testuite");

        // Basic tests of the main functions. All results are expected KO
        `WARNING("Start to launch KO testsuite");
        `CRITICAL("All tests are expected KO");
        `INFO("Test FAIL_IF_NOT");
        `FAIL_IF_NOT(inc);
        @(posedge aclk);
        inc = 1'b1;
        `INFO("Test FAIL_IF");
        `FAIL_IF(inc);
        @(posedge aclk);
        inc = 1'b0;
        `INFO("Test FAIL_IF_NOT");
        `FAIL_IF_NOT(inc);
        `INFO("Test FAIL_IF_EQUAL");
        `FAIL_IF_NOT_EQUAL(out, 8'd0);
        `INFO("Test FAIL_IF_NOT_EQUAL");
        `FAIL_IF_EQUAL(out, 8'd1);

        `ERROR("Test finished");

    `UNIT_TEST_END

    `TEST_SUITE_END

endmodule

